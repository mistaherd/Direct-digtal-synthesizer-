library verilog;
use verilog.vl_types.all;
entity DSS_vlg_check_tst is
    port(
        FSK_OUT         : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end DSS_vlg_check_tst;
