library verilog;
use verilog.vl_types.all;
entity DSS_vlg_vec_tst is
end DSS_vlg_vec_tst;
